module adder(input [31:0] in1, input [31:0] in2, output reg [31:0] adder_out);
	always @ (in1,in2)
	begin
		adder_out=in1+in2;
	end
endmodule

